`include "definitions.vh"

module ALU_control(
    input [1:0] ALUOp,
    input [5:0] funct,
    output reg  [3:0] ALU_control
    );
    always@(*) begin
    
    //your code here
    
    end
endmodule
