`include "definitions.vh"



module ALU(
    input [`WORD-1:0] A,
    input [`WORD-1:0] B,
    input [3:0] ALU_control,
    output reg[`WORD-1:0] ALUresult,
    output zero
    );
    
    assign zero = ;//fill in the blank :)
    
    always@(*) begin
    
    // your code here
    
    end
endmodule
